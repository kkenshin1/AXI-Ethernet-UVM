`ifndef APB_PKG_SVH
`define APB_PKG_SVH

`include "../testbench/apb_agent/apb_transaction.sv"           //APB事务基础结构包

`include "../testbench/apb_agent/apb_master_driver.sv"         //APB MASTER DRIVER
`include "../testbench/apb_agent/apb_master_monitor.sv"        //APB MASTER MONITOR
`include "../testbench/apb_agent/apb_master_sequencer.sv"      //APB MASTER SEQUENCER
`include "../testbench/apb_agent/apb_master_agent.sv"          //APB MASTER AGENT
`include "../testbench/apb_agent/apb_master_seq_lib.sv"        //APB MASTER SEQUENCE LIB

`include "../testbench/apb_agent/apb_reg_adapter.sv"           //APB MASTER REG ADAPTER


`endif
